bplist00�SURL_mfile:///Users/lukehuang/Library/Messages/Attachments/ad/13/BD0AB364-1D40-4646-BE28-B9430808E046/controller.sv                            